library ieee; use ieee.std_logic_1164.all; use ieee.numeric_std.all; entity
icache_ctrl is port( clk, nrst: in std_logic; hit: in std_logic; ramstate: in
std_logic_vector( 1 downto 0); icache_en: out std_logic; memConflict: in std_logic); end icache_ctrl;
architecture instr_cache_ctrl of icache_ctrl is type state_type is(
l1l1l1l1l1l1l1l1l, l1l1l1l1l1l1l1l1l1); signal
ll11l1l11lll1lll11lll11ll1ll1ll1ll11ll11l1ll1111ll11l11111ll111ll11l11ll1ll1l1l111111l1lll1l1ll1l111ll1l1llll11lllll1l1ll11l11ll
,
l1l11l1l111l111lll1l1l1111lllll11111ll11ll1l1l1ll1l1l1111l1l1lll1111ll1ll11llll11llll111l1l11lll111l111111l1lll11l111lllll11lll1
: state_type; begin icache_state: process( clk, nrst) begin if nrst= '0' then
ll11l1l11lll1lll11lll11ll1ll1ll1ll11ll11l1ll1111ll11l11111ll111ll11l11ll1ll1l1l111111l1lll1l1ll1l111ll1l1llll11lllll1l1ll11l11ll
<= l1l1l1l1l1l1l1l1l; elsif rising_edge( clk) then
ll11l1l11lll1lll11lll11ll1ll1ll1ll11ll11l1ll1111ll11l11111ll111ll11l11ll1ll1l1l111111l1lll1l1ll1l111ll1l1llll11lllll1l1ll11l11ll
<=
l1l11l1l111l111lll1l1l1111lllll11111ll11ll1l1l1ll1l1l1111l1l1lll1111ll1ll11llll11llll111l1l11lll111l111111l1lll11l111lllll11lll1
; end if; end process icache_state; nexttstate: process( hit,
ll11l1l11lll1lll11lll11ll1ll1ll1ll11ll11l1ll1111ll11l11111ll111ll11l11ll1ll1l1l111111l1lll1l1ll1l111ll1l1llll11lllll1l1ll11l11ll
, ramstate, memConflict) begin
l1l11l1l111l111lll1l1l1111lllll11111ll11ll1l1l1ll1l1l1111l1l1lll1111ll1ll11llll11llll111l1l11lll111l111111l1lll11l111lllll11lll1
<=
ll11l1l11lll1lll11lll11ll1ll1ll1ll11ll11l1ll1111ll11l11111ll111ll11l11ll1ll1l1l111111l1lll1l1ll1l111ll1l1llll11lllll1l1ll11l11ll
; icache_en <= '0'; case
ll11l1l11lll1lll11lll11ll1ll1ll1ll11ll11l1ll1111ll11l11111ll111ll11l11ll1ll1l1l111111l1lll1l1ll1l111ll1l1llll11lllll1l1ll11l11ll
is when l1l1l1l1l1l1l1l1l => if (hit= '0' and memConflict = '0') then
l1l11l1l111l111lll1l1l1111lllll11111ll11ll1l1l1ll1l1l1111l1l1lll1111ll1ll11llll11llll111l1l11lll111l111111l1lll11l111lllll11lll1
<= l1l1l1l1l1l1l1l1l1; end if; when l1l1l1l1l1l1l1l1l1 => if ramstate /= "01"
then
l1l11l1l111l111lll1l1l1111lllll11111ll11ll1l1l1ll1l1l1111l1l1lll1111ll1ll11llll11llll111l1l11lll111l111111l1lll11l111lllll11lll1
<= l1l1l1l1l1l1l1l1l; icache_en <= '1'; end if; end case; end process
nexttstate; end;
